magic
tech scmos
timestamp 1734090736
<< nwell >>
rect 1175 -15 1191 4
rect 677 -208 705 -180
<< polysilicon >>
rect 1182 -6 1184 -4
rect 1182 -29 1184 -14
rect 1182 -36 1184 -33
rect 686 -190 688 -188
rect 694 -190 696 -188
rect 686 -234 688 -206
rect 694 -213 696 -206
rect 695 -217 696 -213
rect 694 -234 696 -217
rect 686 -240 688 -238
rect 694 -240 696 -238
<< ndiffusion >>
rect 1181 -33 1182 -29
rect 1184 -33 1185 -29
rect 685 -238 686 -234
rect 688 -238 689 -234
rect 693 -238 694 -234
rect 696 -238 697 -234
<< pdiffusion >>
rect 1176 -14 1177 -6
rect 1181 -14 1182 -6
rect 1184 -14 1185 -6
rect 1189 -14 1190 -6
rect 680 -206 681 -190
rect 685 -206 686 -190
rect 688 -206 694 -190
rect 696 -206 697 -190
rect 701 -206 702 -190
<< metal1 >>
rect 540 205 652 211
rect 675 205 689 211
rect -36 184 6 188
rect 617 184 649 188
rect -37 176 1 180
rect 644 176 656 180
rect 638 156 653 162
rect 440 47 444 74
rect 638 47 642 156
rect 685 106 689 205
rect 440 43 586 47
rect 590 43 642 47
rect 655 102 929 106
rect 655 -181 659 102
rect 925 59 929 102
rect 715 38 945 42
rect 1087 19 1157 25
rect 1152 3 1157 19
rect 1152 2 1233 3
rect 857 -2 931 2
rect 1152 -2 1177 2
rect 1181 -2 1185 2
rect 1189 -2 1233 2
rect 1152 -3 1233 -2
rect 1177 -6 1181 -3
rect 1094 -10 1147 -6
rect 1143 -18 1147 -10
rect 1143 -22 1178 -18
rect 1185 -23 1189 -14
rect 1085 -30 1133 -24
rect 1185 -27 1209 -23
rect 1185 -29 1189 -27
rect 1128 -39 1133 -30
rect 1177 -39 1181 -33
rect 1128 -40 1190 -39
rect 1128 -44 1177 -40
rect 1181 -44 1185 -40
rect 1189 -44 1190 -40
rect 1128 -45 1190 -44
rect 729 -51 957 -47
rect 655 -182 704 -181
rect 655 -186 681 -182
rect 685 -186 689 -182
rect 693 -186 697 -182
rect 701 -186 704 -182
rect 655 -187 704 -186
rect 655 -188 659 -187
rect 542 -194 659 -188
rect 681 -190 685 -187
rect 697 -207 701 -206
rect 729 -207 733 -51
rect 697 -210 733 -207
rect -23 -215 19 -211
rect 606 -215 626 -211
rect -9 -223 7 -219
rect 622 -221 626 -215
rect 630 -217 691 -213
rect 701 -221 705 -210
rect 622 -225 682 -221
rect 689 -225 705 -221
rect 689 -234 693 -225
rect 540 -243 556 -237
rect 681 -242 685 -238
rect 697 -242 701 -238
rect 932 -242 938 -66
rect 1052 -210 1058 -62
rect 1205 -103 1209 -27
rect 1228 -80 1233 -3
rect 1228 -86 1276 -80
rect 1205 -107 1250 -103
rect 1403 -122 1521 -120
rect 1403 -126 1558 -122
rect 1516 -128 1558 -126
rect 1198 -147 1250 -143
rect 1446 -149 1488 -145
rect 2075 -149 2125 -145
rect 1446 -151 1450 -149
rect 1411 -155 1450 -151
rect 1459 -165 1463 -153
rect 1440 -169 1463 -165
rect 1143 -196 1248 -192
rect 1052 -216 1260 -210
rect 586 -246 681 -242
rect 685 -246 689 -242
rect 693 -246 697 -242
rect 701 -246 938 -242
rect 1440 -328 1444 -169
rect 2074 -220 2124 -216
rect 1171 -332 1444 -328
rect 1516 -332 1522 -328
rect 1171 -416 1175 -332
rect -5 -420 1175 -416
rect 544 -601 603 -595
rect -18 -622 24 -618
rect 619 -622 857 -618
rect -9 -630 3 -626
rect 546 -732 560 -731
rect 546 -736 556 -732
rect 546 -737 560 -736
rect 541 -1012 603 -1006
rect -22 -1033 20 -1029
rect 614 -1033 1202 -1029
rect -9 -1041 3 -1037
rect 544 -1148 550 -1142
<< metal2 >>
rect -9 -219 -5 176
rect 586 -199 590 43
rect 599 -189 603 -188
rect 586 -203 595 -199
rect -9 -416 -5 -223
rect 590 -231 595 -203
rect 586 -236 595 -231
rect 586 -237 590 -236
rect 552 -238 590 -237
rect 556 -242 590 -238
rect 552 -243 586 -242
rect -9 -626 -5 -420
rect -9 -1037 -5 -630
rect 586 -731 590 -246
rect 556 -732 590 -731
rect 560 -736 590 -732
rect 556 -737 590 -736
rect 586 -1020 590 -737
rect 599 -596 603 -193
rect 630 -213 634 184
rect 673 176 715 180
rect 644 -221 648 176
rect 711 42 715 176
rect 599 -1007 603 -600
rect 853 -618 857 -2
rect 1143 -192 1147 -22
rect 599 -1012 603 -1011
rect 586 -1024 597 -1020
rect 593 -1040 597 -1024
rect 1198 -1029 1202 -147
rect 1338 -318 1344 -210
rect 1338 -323 1457 -318
rect 1452 -328 1457 -323
rect 1452 -332 1516 -328
rect 586 -1044 597 -1040
rect 586 -1142 590 -1044
rect 544 -1143 590 -1142
rect 544 -1147 545 -1143
rect 549 -1147 590 -1143
rect 544 -1148 590 -1147
<< ntransistor >>
rect 1182 -33 1184 -29
rect 686 -238 688 -234
rect 694 -238 696 -234
<< ptransistor >>
rect 1182 -14 1184 -6
rect 686 -206 688 -190
rect 694 -206 696 -190
<< polycontact >>
rect 1178 -22 1182 -18
rect 682 -225 686 -221
rect 691 -217 695 -213
<< ndcontact >>
rect 1177 -33 1181 -29
rect 1185 -33 1189 -29
rect 681 -238 685 -234
rect 689 -238 693 -234
rect 697 -238 701 -234
<< pdcontact >>
rect 1177 -14 1181 -6
rect 1185 -14 1189 -6
rect 681 -206 685 -190
rect 697 -206 701 -190
<< m2contact >>
rect 586 43 590 47
rect 711 38 715 42
rect 853 -2 857 2
rect -9 -420 -5 -416
rect 556 -736 560 -732
<< psubstratepcontact >>
rect 1177 -44 1181 -40
rect 1185 -44 1189 -40
rect 681 -246 685 -242
rect 689 -246 693 -242
rect 697 -246 701 -242
<< highvoltnsubcontact >>
rect 1177 -2 1181 2
rect 1185 -2 1189 2
rect 681 -186 685 -182
rect 689 -186 693 -182
rect 697 -186 701 -182
<< pad >>
rect 630 184 634 188
rect -9 176 -5 180
rect 599 -193 603 -189
rect -9 -223 -5 -219
rect 552 -242 556 -238
rect -9 -630 -5 -626
rect 586 -246 590 -242
rect 630 -217 634 -213
rect 644 176 648 180
rect 644 -225 648 -221
rect 599 -600 603 -596
rect 1143 -22 1147 -18
rect 1143 -196 1147 -192
rect 1198 -147 1202 -143
rect 853 -622 857 -618
rect 599 -1011 603 -1007
rect -9 -1041 -5 -1037
rect 1516 -332 1522 -328
rect 1198 -1033 1202 -1029
rect 545 -1147 549 -1143
use dff dff_0
timestamp 1734089879
transform 1 0 29 0 1 57
box -29 -57 588 155
use nand nand_0
timestamp 1731253790
transform 1 0 662 0 1 192
box -16 -36 15 20
use mux mux_0
timestamp 1734027179
transform 1 0 984 0 1 10
box -55 -81 110 56
use dff dff_1
timestamp 1734089879
transform 1 0 30 0 1 -342
box -29 -57 588 155
use mux mux_1
timestamp 1734027179
transform 1 0 1301 0 1 -135
box -55 -81 110 56
use dff dff_4
timestamp 1734089879
transform 1 0 1488 0 1 -276
box -29 -57 588 155
use dff dff_2
timestamp 1734089879
transform 1 0 32 0 1 -749
box -29 -57 588 155
use dff dff_3
timestamp 1734089879
transform 1 0 30 0 1 -1160
box -29 -57 588 155
<< labels >>
rlabel metal1 2115 -218 2115 -218 1 Qnot
rlabel metal1 2114 -147 2114 -147 1 r_result
rlabel metal1 1438 -153 1438 -153 1 node9
rlabel metal2 1200 -420 1200 -420 1 node8
rlabel metal1 1207 -87 1207 -87 1 node7
rlabel metal1 1137 -8 1137 -8 1 node6
rlabel metal2 855 -377 855 -377 1 node5
rlabel metal1 784 -49 784 -49 1 node4
rlabel metal1 789 40 789 40 1 node3
rlabel metal1 676 -244 676 -244 1 gnd
rlabel metal1 669 -184 669 -184 1 vdd
rlabel metal1 632 186 632 186 1 node1
rlabel metal1 -31 178 -31 178 1 clk
rlabel metal1 -31 186 -31 186 3 input_a
rlabel metal1 -18 -213 -18 -213 1 input_b
rlabel metal1 -17 -1031 -17 -1031 1 ins_1
rlabel metal1 -15 -620 -15 -620 1 ins_0
rlabel pad 646 -223 646 -223 1 node2
<< end >>
