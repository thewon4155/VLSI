magic
tech scmos
timestamp 1731253790
<< nwell >>
rect -13 1 15 20
<< polysilicon >>
rect -4 10 -2 12
rect 4 10 6 12
rect -4 -23 -2 2
rect 4 -12 6 2
rect 4 -23 6 -16
rect -4 -29 -2 -27
rect 4 -29 6 -27
<< ndiffusion >>
rect -5 -27 -4 -23
rect -2 -27 -1 -23
rect 3 -27 4 -23
rect 6 -27 7 -23
<< pdiffusion >>
rect -10 2 -9 10
rect -5 2 -4 10
rect -2 2 -1 10
rect 3 2 4 10
rect 6 2 7 10
rect 11 2 12 10
<< metal1 >>
rect -12 18 14 19
rect -12 14 -9 18
rect -5 14 -1 18
rect 3 14 7 18
rect 11 14 14 18
rect -12 13 14 14
rect -9 10 -5 13
rect 7 10 11 13
rect -1 -4 3 2
rect -16 -8 -8 -4
rect -16 -16 4 -12
rect 11 -27 15 -16
rect -9 -30 -5 -27
rect -10 -31 12 -30
rect -10 -35 -9 -31
rect -5 -35 -1 -31
rect 3 -35 7 -31
rect 11 -35 12 -31
rect -10 -36 12 -35
<< metal2 >>
rect 3 -4 11 0
rect 11 -12 15 -4
<< ntransistor >>
rect -4 -27 -2 -23
rect 4 -27 6 -23
<< ptransistor >>
rect -4 2 -2 10
rect 4 2 6 10
<< polycontact >>
rect -8 -8 -4 -4
rect 4 -16 8 -12
<< ndcontact >>
rect -9 -27 -5 -23
rect -1 -27 3 -23
rect 7 -27 11 -23
<< pdcontact >>
rect -9 2 -5 10
rect -1 2 3 10
rect 7 2 11 10
<< m2contact >>
rect 11 -16 15 -12
<< psubstratepcontact >>
rect -9 -35 -5 -31
rect -1 -35 3 -31
rect 7 -35 11 -31
<< highvoltnsubcontact >>
rect -9 14 -5 18
rect -1 14 3 18
rect 7 14 11 18
<< pad >>
rect -1 -4 3 0
rect 11 -4 15 0
<< labels >>
rlabel metal1 5 16 5 16 5 vdd
rlabel metal1 5 -33 5 -33 1 gnd
rlabel metal1 -10 -6 -10 -6 1 in1
rlabel metal1 -9 -14 -9 -14 1 in2
rlabel metal2 13 -9 13 -9 7 out
<< end >>
