magic
tech scmos
timestamp 1731503720
<< nwell >>
rect -108 -81 -82 -61
<< polysilicon >>
rect -85 6 -65 10
rect -130 -2 -108 2
rect -85 -2 -66 2
rect -131 -17 -104 -16
rect -131 -21 -130 -17
rect -126 -21 -109 -17
rect -105 -21 -104 -17
rect -131 -22 -104 -21
rect -77 -28 -73 -11
rect -62 -26 -58 -13
rect -8 -17 15 -16
rect -8 -21 -7 -17
rect -3 -21 10 -17
rect 14 -21 15 -17
rect -8 -22 15 -21
rect -62 -65 -58 -49
rect 60 -65 79 -61
rect -96 -72 -94 -70
rect -96 -92 -94 -80
rect -96 -98 -94 -96
rect -8 -104 19 -103
rect -8 -108 -7 -104
rect -3 -108 14 -104
rect 18 -108 19 -104
rect -8 -109 19 -108
<< ndiffusion >>
rect -97 -96 -96 -92
rect -94 -96 -93 -92
<< pdiffusion >>
rect -103 -80 -101 -72
rect -97 -80 -96 -72
rect -94 -80 -93 -72
rect -89 -80 -87 -72
<< metal1 >>
rect -77 27 -46 33
rect -20 27 18 33
rect -144 6 -89 10
rect -144 -2 -134 2
rect -137 -17 -125 -16
rect -137 -21 -130 -17
rect -126 -21 -125 -17
rect -137 -22 -125 -21
rect -137 -100 -131 -22
rect -121 -84 -117 6
rect -104 -2 -89 2
rect -77 -7 -73 27
rect -61 6 -50 10
rect -23 6 14 10
rect 41 6 98 10
rect -62 -2 -50 2
rect 2 -2 17 2
rect -62 -9 -58 -2
rect -110 -17 -44 -16
rect -110 -21 -109 -17
rect -105 -19 -44 -17
rect -22 -17 -3 -16
rect -22 -19 -7 -17
rect -105 -21 -7 -19
rect -110 -22 -3 -21
rect -77 -54 -73 -32
rect -62 -45 -58 -30
rect 2 -30 6 -2
rect 10 -17 20 -16
rect 14 -21 20 -17
rect 10 -22 20 -21
rect 2 -34 60 -30
rect -77 -60 -45 -54
rect -19 -60 22 -54
rect -77 -63 -73 -60
rect -103 -64 -73 -63
rect -103 -68 -101 -64
rect -97 -68 -93 -64
rect -89 -68 -73 -64
rect 56 -61 60 -34
rect -103 -69 -73 -68
rect -101 -72 -97 -69
rect -121 -88 -100 -84
rect -93 -85 -89 -80
rect -62 -77 -58 -69
rect -62 -81 -48 -77
rect -22 -81 19 -77
rect 56 -85 60 -65
rect -93 -89 -49 -85
rect 4 -89 18 -85
rect 45 -89 60 -85
rect -93 -92 -89 -89
rect -101 -100 -97 -96
rect -137 -101 -62 -100
rect -137 -105 -101 -101
rect -97 -105 -93 -101
rect -89 -103 -62 -101
rect -89 -105 -42 -103
rect -137 -106 -42 -105
rect -66 -109 -42 -106
rect -21 -104 -3 -103
rect -21 -108 -7 -104
rect -21 -109 -3 -108
rect 4 -117 8 -89
rect 14 -104 24 -103
rect 18 -108 24 -104
rect 14 -109 24 -108
rect 67 -117 71 6
rect 83 -65 99 -61
rect 4 -121 71 -117
<< ntransistor >>
rect -96 -96 -94 -92
<< ptransistor >>
rect -96 -80 -94 -72
<< polycontact >>
rect -89 6 -85 10
rect -65 6 -61 10
rect -134 -2 -130 2
rect -108 -2 -104 2
rect -89 -2 -85 2
rect -66 -2 -62 2
rect -77 -11 -73 -7
rect -130 -21 -126 -17
rect -109 -21 -105 -17
rect -77 -32 -73 -28
rect -62 -13 -58 -9
rect -7 -21 -3 -17
rect 10 -21 14 -17
rect -62 -30 -58 -26
rect -62 -49 -58 -45
rect 56 -65 60 -61
rect 79 -65 83 -61
rect -62 -69 -58 -65
rect -100 -88 -96 -84
rect -7 -108 -3 -104
rect 14 -108 18 -104
<< ndcontact >>
rect -101 -96 -97 -92
rect -93 -96 -89 -92
<< pdcontact >>
rect -101 -80 -97 -72
rect -93 -80 -89 -72
<< psubstratepcontact >>
rect -101 -105 -97 -101
rect -93 -105 -89 -101
<< highvoltnsubcontact >>
rect -101 -68 -97 -64
rect -93 -68 -89 -64
<< pad >>
rect -23 6 -19 10
rect 41 6 45 10
rect -22 -81 -18 -77
use nand nand_0
timestamp 1731253790
transform 1 0 -34 0 1 14
box -16 -36 15 20
use nand nand_1
timestamp 1731253790
transform 1 0 30 0 1 14
box -16 -36 15 20
use nand nand_2
timestamp 1731253790
transform 1 0 -33 0 1 -73
box -16 -36 15 20
use nand nand_3
timestamp 1731253790
transform 1 0 34 0 1 -73
box -16 -36 15 20
<< labels >>
rlabel metal1 -95 -66 -95 -66 1 vdd
rlabel metal1 -95 -103 -95 -103 1 gnd
rlabel metal1 -142 8 -142 8 3 input1
rlabel metal1 -142 0 -142 0 3 input2
rlabel metal1 91 8 91 8 1 Q
rlabel metal1 93 -63 93 -63 1 Qnot
rlabel metal1 1 8 1 8 1 node1
rlabel metal1 3 -79 3 -79 1 node2
rlabel metal1 -65 -87 -65 -87 1 node3
<< end >>
