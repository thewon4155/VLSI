magic
tech scmos
timestamp 1731503720
<< nwell >>
rect -43 -39 -21 -19
<< polysilicon >>
rect -23 28 0 32
rect -64 20 -51 24
rect -23 20 -4 24
rect -4 -19 0 -1
rect 97 -28 116 -24
rect -33 -30 -31 -28
rect -33 -50 -31 -38
rect -33 -57 -31 -54
<< ndiffusion >>
rect -34 -54 -33 -50
rect -31 -54 -30 -50
<< pdiffusion >>
rect -39 -38 -38 -30
rect -34 -38 -33 -30
rect -31 -38 -30 -30
rect -26 -38 -25 -30
<< metal1 >>
rect -16 49 4 55
rect 29 49 55 55
rect -77 28 -27 32
rect -77 20 -68 24
rect -60 -43 -56 28
rect -47 20 -27 24
rect -16 -9 -11 49
rect 4 28 7 32
rect 31 28 51 32
rect 78 30 131 34
rect -4 3 0 20
rect 37 20 61 24
rect 37 -5 42 20
rect -16 -15 4 -9
rect 30 -15 34 -9
rect 37 -10 97 -5
rect -16 -20 -11 -15
rect -41 -21 -11 -20
rect -41 -25 -38 -21
rect -34 -25 -30 -21
rect -26 -25 -11 -21
rect -41 -26 -11 -25
rect 30 -21 59 -15
rect -38 -30 -34 -26
rect -4 -32 0 -23
rect 92 -24 97 -10
rect -4 -36 8 -32
rect 27 -36 47 -32
rect 92 -35 97 -28
rect -30 -40 -26 -38
rect 43 -38 47 -36
rect -60 -47 -37 -43
rect -30 -44 0 -40
rect 43 -42 61 -38
rect 80 -39 97 -35
rect -30 -50 -26 -44
rect 43 -50 54 -46
rect -38 -58 -34 -54
rect -40 -59 -24 -58
rect -40 -63 -38 -59
rect -34 -63 -30 -59
rect -26 -63 -24 -59
rect -40 -64 -24 -63
rect 43 -76 47 -50
rect 105 -76 110 30
rect 121 -28 132 -24
rect 43 -80 110 -76
<< ntransistor >>
rect -33 -54 -31 -50
<< ptransistor >>
rect -33 -38 -31 -30
<< polycontact >>
rect -27 28 -23 32
rect 0 28 4 32
rect -68 20 -64 24
rect -51 20 -47 24
rect -27 20 -23 24
rect -4 20 0 24
rect -4 -1 0 3
rect -4 -23 0 -19
rect 92 -28 97 -24
rect 116 -28 121 -24
rect -37 -47 -33 -43
<< ndcontact >>
rect -38 -54 -34 -50
rect -30 -54 -26 -50
<< pdcontact >>
rect -38 -38 -34 -30
rect -30 -38 -26 -30
<< m2contact >>
rect 27 28 31 32
<< psubstratepcontact >>
rect -38 -63 -34 -59
rect -30 -63 -26 -59
<< highvoltnsubcontact >>
rect -38 -25 -34 -21
rect -30 -25 -26 -21
<< pad >>
rect 78 30 82 33
rect 27 -36 31 -32
rect 80 -39 84 -35
use nand nand_0
timestamp 1731253790
transform 1 0 16 0 1 36
box -16 -36 15 20
use nand nand_2
timestamp 1731253790
transform 1 0 67 0 1 36
box -16 -36 15 20
use nand nand_1
timestamp 1731253790
transform 1 0 16 0 1 -28
box -16 -36 15 20
use nand nand_3
timestamp 1731253790
transform 1 0 69 0 1 -34
box -16 -36 15 20
<< labels >>
rlabel metal1 44 52 44 52 5 Vdd
rlabel metal1 -32 -62 -32 -62 1 gnd
rlabel metal1 -76 30 -76 30 3 D
rlabel metal1 -76 22 -76 22 3 CLK
rlabel metal1 46 30 46 30 1 node1
rlabel metal1 43 -35 43 -35 1 node2
rlabel metal1 -9 -41 -9 -41 1 node3
rlabel metal1 109 31 109 31 1 Q
rlabel metal1 127 -26 127 -26 7 Qnot
<< end >>
